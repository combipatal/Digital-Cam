// Digital camera implementation #4
// Features:
// > Normal video mode
// > Realtime edge detection video mode

module digital_cam_impl4(
    input clk_50,
    input btn_RESET, // KEY0; manual reset
    input slide_sw_resend_reg_values, // rewrite all OV7670's registers
    input slide_sw_NORMAL_OR_EDGEDETECT, // 0 normal, 1 edge detection

    output vga_hsync,
    output vga_vsync,
    output [7:0] vga_r,
    output [7:0] vga_g,
    output [7:0] vga_b,
    output vga_blank_N,
    output vga_sync_N,
    output vga_CLK,

    input ov7670_pclk,
    output ov7670_xclk,
    input ov7670_vsync,
    input ov7670_href,
    input [7:0] ov7670_data,
    output ov7670_sioc,
    inout ov7670_siod,
    output ov7670_pwdn,
    output ov7670_reset,

    output LED_config_finished, // lets us know camera registers are now written
    output LED_dll_locked, // PLL is locked now
    output LED_done
);

    // PLL outputs
    wire clk_100;       // c0: 100 MHz
    wire clk_100_3ns;   // c1: 100 MHz with phase adjustment of -3ns
    wire clk_50_camera; // c2: 50 MHz
    wire clk_25_vga;    // c3: 25 MHz
    wire dll_locked;

    // Signals that need to be assigned in always blocks
    reg done_BW_reg = 1'b0;
    reg done_ED_reg = 1'b0;
    reg done_capture_new_frame_reg = 1'b0;
    wire done_BW_from_module;
    wire done_ED_from_module;
    wire done_capture_new_frame_from_module;

    // Connect module outputs to internal registers
    always @(posedge clk_25_vga) begin
        done_BW_reg <= done_BW_from_module;
        done_ED_reg <= done_ED_from_module;
        done_capture_new_frame_reg <= done_capture_new_frame_from_module;
    end

    // Buffer 1 signals
    reg wren_buf_1 = 1'b0;
    reg [16:0] wraddress_buf_1 = 17'b0;
    reg [11:0] wrdata_buf_1 = 12'b0;
    reg [16:0] rdaddress_buf_1 = 17'b0;
    wire [11:0] rddata_buf_1;

    // Signals generated by different entities will be multiplexed into the
    // inputs above of buffer 1
    wire [16:0] rdaddress_buf12_from_addr_gen; // muxed to both buf1 and buf2
    wire [16:0] rdaddress_buf1_from_do_BW;
    wire [16:0] rdaddress_buf1_from_do_ED;
    wire wren_buf1_from_ov7670_capture;
    wire [16:0] wraddress_buf1_from_ov7670_capture;
    wire [11:0] wrdata_buf1_from_ov7670_capture;
    wire wren_buf1_from_do_BW;
    wire [16:0] wraddress_buf1_from_do_BW;
    wire [11:0] wrdata_buf1_from_do_BW;

    // Buffer 2 signals
    reg wren_buf_2 = 1'b0;
    reg [16:0] wraddress_buf_2 = 17'b0;
    reg [11:0] wrdata_buf_2 = 12'b0;
    reg [16:0] rdaddress_buf_2 = 17'b0;
    wire [11:0] rddata_buf_2;

    // Signals generated by different entities will be multiplexed into the
    // inputs above of buffer 2
    // Signals to control buffer 2 when reading it, do edge detection, and then write back into it
    wire wren_buf2_from_do_ED;
    wire [16:0] wraddress_buf2_from_do_ED;
    wire [11:0] wrdata_buf2_from_do_ED;

    // User controls
    wire resend_reg_values;
    wire normal_or_edgedetect;
    wire reset_manual; // by user via KEY0 push button
    reg reset_automatic = 1'b0; // TODO: make it 1 for 2 clock cycles, then permanently to 0
    wire reset_global; // combination of previous two
    reg reset_BW_entity = 1'b0;
    reg reset_ED_entity = 1'b0;

    reg call_black_white = 1'b0;
    reg call_edge_detection = 1'b0;
    reg call_black_white_synchronized = 1'b0;
    reg call_edge_detection_synchronized = 1'b0;

    // RGB related
    wire [7:0] red, green, blue;
    wire activeArea;
    wire nBlank;
    wire vSync;
    // data_to_rgb should the multiplexing of rddata_buf_1 (when displaying
    // video directly) or rddata_buf_2 (for realtime edge detection video mode)
    reg [11:0] data_to_rgb = 12'b0;

    // Top level control
    localparam [2:0]
        S0_RESET = 3'b000,
        S1_RESET_BW = 3'b001,
        S2_PROCESS_BW = 3'b010,
        S3_DONE_BW = 3'b011,
        S4_RESET_ED = 3'b100,
        S5_PROCESS_ED = 3'b101,
        S6_DONE_ED = 3'b110,
        S7_NORMAL_VIDEO_MODE = 3'b111;

    reg [2:0] state_current = S0_RESET, state_next;

    // State register; process #1
    always @(posedge clk_25_vga, posedge reset_global) begin
        if (reset_global) begin
            state_current <= S0_RESET;
        end else begin
            state_current <= state_next;
        end
    end

    // Next state and output logic; process #2
    always @* begin
        state_next = state_current;
        reset_BW_entity = 1'b0;
        reset_ED_entity = 1'b0;
        call_black_white = 1'b0;
        call_edge_detection = 1'b0;

        case (state_current)
            S0_RESET: begin
                reset_BW_entity = 1'b1;
                reset_ED_entity = 1'b1;
                if (normal_or_edgedetect == 1'b0) begin // normal video mode
                    state_next = S7_NORMAL_VIDEO_MODE;
                    data_to_rgb = rddata_buf_1; // show buf1 on VGA monitor
                    // signals of buf1
                    wren_buf_1 = wren_buf1_from_ov7670_capture;
                    wraddress_buf_1 = wraddress_buf1_from_ov7670_capture;
                    wrdata_buf_1 = wrdata_buf1_from_ov7670_capture;
                    rdaddress_buf_1 = rdaddress_buf12_from_addr_gen;
                    // signals of buf2
                    wren_buf_2 = 1'b0; // disabled
                    wraddress_buf_2 = wraddress_buf2_from_do_ED; // don't care
                    wrdata_buf_2 = wrdata_buf2_from_do_ED; // don't care
                    rdaddress_buf_2 = rdaddress_buf12_from_addr_gen;
                end else begin // realtime edge detection video mode
                    state_next = S1_RESET_BW;
                    data_to_rgb = rddata_buf_2; // show buf2 on VGA monitor
                    // signals of buf1
                    wren_buf_1 = wren_buf1_from_do_BW;
                    wraddress_buf_1 = wraddress_buf1_from_do_BW;
                    wrdata_buf_1 = wrdata_buf1_from_do_BW;
                    rdaddress_buf_1 = rdaddress_buf1_from_do_BW;
                    // signals of buf2
                    wren_buf_2 = 1'b0; // disabled
                    wraddress_buf_2 = wraddress_buf2_from_do_ED; // don't care
                    wrdata_buf_2 = wrdata_buf2_from_do_ED; // don't care
                    rdaddress_buf_2 = rdaddress_buf12_from_addr_gen;
                end
            end

            // Next states, except the last one, are went thru only during realtime
            // edge detection video mode
            S1_RESET_BW: begin
                reset_BW_entity = 1'b1;
                state_next = S2_PROCESS_BW;
                data_to_rgb = rddata_buf_2; // show buf2 on VGA monitor
                // signals of buf1
                wren_buf_1 = wren_buf1_from_do_BW;
                wraddress_buf_1 = wraddress_buf1_from_do_BW;
                wrdata_buf_1 = wrdata_buf1_from_do_BW;
                rdaddress_buf_1 = rdaddress_buf1_from_do_BW;
                // signals of buf2
                wren_buf_2 = 1'b0; // disabled
                wraddress_buf_2 = wraddress_buf2_from_do_ED; // don't care
                wrdata_buf_2 = wrdata_buf2_from_do_ED; // don't care
                rdaddress_buf_2 = rdaddress_buf12_from_addr_gen;
            end

            S2_PROCESS_BW: begin
                call_black_white = 1'b1; // used to generate call_black_white_synchronized
                if (done_BW_reg == 1'b0) begin
                    state_next = S2_PROCESS_BW;
                end else begin
                    state_next = S3_DONE_BW;
                end
                data_to_rgb = rddata_buf_2; // show buf2 on VGA monitor
                // signals of buf1
                wren_buf_1 = wren_buf1_from_do_BW;
                wraddress_buf_1 = wraddress_buf1_from_do_BW;
                wrdata_buf_1 = wrdata_buf1_from_do_BW;
                rdaddress_buf_1 = rdaddress_buf1_from_do_BW;
                // signals of buf2
                wren_buf_2 = 1'b0; // disabled
                wraddress_buf_2 = wraddress_buf2_from_do_ED; // don't care
                wrdata_buf_2 = wrdata_buf2_from_do_ED; // don't care
                rdaddress_buf_2 = rdaddress_buf12_from_addr_gen;
            end

            S3_DONE_BW: begin
                reset_BW_entity = 1'b1; // to put it in idle immediately; done BW is thus just one cycle
                state_next = S4_RESET_ED;
                data_to_rgb = rddata_buf_2; // show buf2 on VGA monitor
                // signals of buf1
                wren_buf_1 = 1'b0; // disabled
                wraddress_buf_1 = wraddress_buf1_from_do_BW;
                wrdata_buf_1 = wrdata_buf1_from_do_BW;
                rdaddress_buf_1 = rdaddress_buf1_from_do_BW;
                // signals of buf2
                wren_buf_2 = 1'b0; // disabled
                wraddress_buf_2 = wraddress_buf2_from_do_ED; // don't care
                wrdata_buf_2 = wrdata_buf2_from_do_ED; // don't care
                rdaddress_buf_2 = rdaddress_buf12_from_addr_gen;
            end

            S4_RESET_ED: begin
                reset_ED_entity = 1'b1;
                state_next = S5_PROCESS_ED;
                data_to_rgb = rddata_buf_2; // show buf2 on VGA monitor
                // signals of buf1
                wren_buf_1 = 1'b0; // disabled
                wraddress_buf_1 = wraddress_buf1_from_do_BW; // don't care
                wrdata_buf_1 = wrdata_buf1_from_do_BW; // don't care
                rdaddress_buf_1 = rdaddress_buf1_from_do_ED; // here we start reading from buf1
                // signals of buf2
                wren_buf_2 = wren_buf2_from_do_ED;
                wraddress_buf_2 = wraddress_buf2_from_do_ED;
                wrdata_buf_2 = wrdata_buf2_from_do_ED;
                rdaddress_buf_2 = rdaddress_buf12_from_addr_gen;
            end

            S5_PROCESS_ED: begin
                call_edge_detection = 1'b1;
                if (done_ED_reg == 1'b0) begin
                    state_next = S5_PROCESS_ED;
                end else begin
                    state_next = S6_DONE_ED;
                end
                data_to_rgb = rddata_buf_2; // show buf2 on VGA monitor
                // signals of buf1
                wren_buf_1 = 1'b0; // disabled
                wraddress_buf_1 = wraddress_buf1_from_do_BW; // don't care
                wrdata_buf_1 = wrdata_buf1_from_do_BW; // don't care
                rdaddress_buf_1 = rdaddress_buf1_from_do_ED;
                // signals of buf2
                wren_buf_2 = wren_buf2_from_do_ED;
                wraddress_buf_2 = wraddress_buf2_from_do_ED;
                wrdata_buf_2 = wrdata_buf2_from_do_ED;
                rdaddress_buf_2 = rdaddress_buf12_from_addr_gen;
            end

            S6_DONE_ED: begin
                reset_ED_entity = 1'b1; // to put it in idle immediately; done ED is thus just one cycle
                state_next = S7_NORMAL_VIDEO_MODE; // S0_RESET;
                data_to_rgb = rddata_buf_2; // show buf2 on VGA monitor
                // signals of buf1
                wren_buf_1 = 1'b0; // disabled
                wraddress_buf_1 = wraddress_buf1_from_do_BW; // don't care
                wrdata_buf_1 = wrdata_buf1_from_do_BW; // don't care
                rdaddress_buf_1 = rdaddress_buf12_from_addr_gen;
                // signals of buf2
                wren_buf_2 = 1'b0; // disabled
                wraddress_buf_2 = wraddress_buf2_from_do_ED;
                wrdata_buf_2 = wrdata_buf2_from_do_ED;
                rdaddress_buf_2 = rdaddress_buf12_from_addr_gen;
            end

            // At this moment, we are done with one sequence of BW+ED; so, now
            // allow a new frame from camera module into buf1
            S7_NORMAL_VIDEO_MODE: begin
                if (normal_or_edgedetect == 1'b0) begin // normal video mode
                    state_next = S7_NORMAL_VIDEO_MODE;
                    data_to_rgb = rddata_buf_1; // show buf1 on VGA monitor
                    // signals of buf1
                    wren_buf_1 = wren_buf1_from_ov7670_capture;
                    wraddress_buf_1 = wraddress_buf1_from_ov7670_capture;
                    wrdata_buf_1 = wrdata_buf1_from_ov7670_capture;
                    rdaddress_buf_1 = rdaddress_buf12_from_addr_gen;
                    // signals of buf2
                    wren_buf_2 = 1'b0; // disabled
                    wraddress_buf_2 = wraddress_buf2_from_do_ED; // don't care
                    wrdata_buf_2 = wrdata_buf2_from_do_ED; // don't care
                    rdaddress_buf_2 = rdaddress_buf12_from_addr_gen;
                end else begin // realtime edge detection video mode
                    if (done_capture_new_frame_reg == 1'b0) begin
                        state_next = S7_NORMAL_VIDEO_MODE; // stay here till we get a complete frame from camera
                    end else begin
                        state_next = S0_RESET;
                    end
                    data_to_rgb = rddata_buf_2; // show buf2 on VGA monitor
                    // signals of buf1
                    wren_buf_1 = wren_buf1_from_ov7670_capture;
                    wraddress_buf_1 = wraddress_buf1_from_ov7670_capture;
                    wrdata_buf_1 = wrdata_buf1_from_ov7670_capture;
                    rdaddress_buf_1 = rdaddress_buf12_from_addr_gen;
                    // signals of buf2
                    wren_buf_2 = 1'b0; // disabled
                    wraddress_buf_2 = wraddress_buf2_from_do_ED; // don't care
                    wrdata_buf_2 = wrdata_buf2_from_do_ED; // don't care
                    rdaddress_buf_2 = rdaddress_buf12_from_addr_gen;
                end
            end

            default: begin
                state_next = S0_RESET;
            end
        endcase
    end

    // LEDs; LED_config_finished is driven directly by entity ov7670_controller
    assign LED_dll_locked = reset_global; // LEDRed[0] notifies user
    assign LED_done = (done_BW | done_ED); // output of top-level entity

    // Clocks generation
    my_altpll four_clocks_pll(
        .areset(1'b0), // reset_general?
        .inclk0(clk_50),
        .c0(clk_100),
        .c1(clk_100_3ns), // not needed anymore
        .c2(clk_50_camera),
        .c3(clk_25_vga),
        .locked(dll_locked) // drives an LED and SDRAM controller
    );

    // Debouncing slide switches, to get clean signals
    debounce debounce_resend(
        .clk(clk_100),
        .reset(reset_global),
        .sw(slide_sw_resend_reg_values),
        .db(resend_reg_values)
    );

    debounce debounce_normal_or_edgedetect(
        .clk(clk_100),
        .reset(reset_global),
        .sw(slide_sw_NORMAL_OR_EDGEDETECT),
        .db(normal_or_edgedetect) // 0 is normal video video; 1 is edge detection in video mode
    );

    // Take the inverted push button because KEY0 on DE2-115 board generates
    // a signal 111000111; with 1 with not pressed and 0 when pressed/pushed
    assign reset_manual = ~btn_RESET; // KEY0
    // First thing when the system is powered on, I should automatically
    // reset everything for a few clock cycles
    assign reset_global = (reset_manual | reset_automatic);

    // Video frames are buffered into buf1; from here, a frame is taken
    // and applied BW on it; written back into buf1; then, as second phase
    // buf1 is read from by ED, which places result into buf2; from where
    // it is displayed on VGA monitor; in normal video mode the above is not
    // done; buf1 is displayed directly on VGA monitor instead
    // VERY IMPORTANT NOTE:
    // initially, in implementations 1-3, I had "wrclock => ov7670_pclk,"
    // because the only entity to write into buf1 was camera module; here, however
    // BW also write its result; so, I could have either "muxed" ov7670_pclk AND clk_25_vga
    // to feed "wrclock", or, just use directly clk_25_vga, which happens to be the same
    // as ov7670_pclk in this particular instance
    frame_buffer frame_buf_1(
        .rdaddress(rdaddress_buf_1),
        .rdclock(clk_25_vga),
        .q(rddata_buf_1), // goes to data_to_rgb thru mux
        .wrclock(clk_25_vga), // ov7670_pclk, clock from camera module
        .wraddress(wraddress_buf_1),
        .data(wrdata_buf_1),
        .wren(wren_buf_1)
    );

    // Buf2 is used to store result of ED, which read from buf1
    frame_buffer frame_buf_2(
        .rdaddress(rdaddress_buf_2),
        .rdclock(clk_25_vga),
        .q(rddata_buf_2), // goes to data_to_rgb thru mux
        .wrclock(clk_25_vga),
        .wraddress(wraddress_buf_2),
        .data(wrdata_buf_2),
        .wren(wren_buf_2)
    );

    // Camera module related blocks
    ov7670_controller ov7670_controller_inst(
        .clk(clk_50_camera),
        .resend(resend_reg_values), // debounced
        .config_finished(LED_config_finished), // LEDRed[1] notifies user
        .sioc(ov7670_sioc),
        .siod(ov7670_siod),
        .reset(ov7670_reset),
        .pwdn(ov7670_pwdn),
        .xclk(ov7670_xclk)
    );

    ov7670_capture ov7670_capture_inst(
        .pclk(ov7670_pclk),
        .vsync(ov7670_vsync),
        .href(ov7670_href),
        .d(ov7670_data),
        .addr(wraddress_buf1_from_ov7670_capture), // wraddress_buf_1 driven by ov7670_capture
        .dout(wrdata_buf1_from_ov7670_capture), // wrdata_buf_1 driven by ov7670_capture
        .we(wren_buf1_from_ov7670_capture), // goes to mux of wren_buf_1
        .end_of_frame(done_capture_new_frame_from_module) // new out signal; did not have it before
    );

    // VGA related stuff
    VGA VGA_inst(
        .CLK25(clk_25_vga),
        .clkout(vga_CLK),
        .Hsync(vga_hsync),
        .Vsync(vsync),
        .Nblank(nBlank),
        .Nsync(vga_sync_N),
        .activeArea(activeArea)
    );

    RGB RGB_inst(
        .Din(data_to_rgb), // comes from either rddata_buf_1 or rddata_buf_2
        .Nblank(activeArea),
        .R(red),
        .G(green),
        .B(blue)
    );

    // VGA related signals
    assign vga_r = red[7:0];
    assign vga_g = green[7:0];
    assign vga_b = blue[7:0];
    assign vga_vsync = vsync;
    assign vga_blank_N = nBlank;

    // "General purpose" address generator
    Address_Generator Address_Generator_inst(
        .rst_i(1'b0),
        .CLK25(clk_25_vga),
        .enable(activeArea),
        .vsync(vsync),
        .address(rdaddress_buf12_from_addr_gen) // goes to muxes of rdaddress_buf_1 and rdaddress_buf_2
    );

    // Generate pulse signals only when vsync is '0' to take a frame from a given buffer
    // synchronized with the beginning of it; otherwise, pixels may be picked-up
    // from different frames
    always @* begin
        call_black_white_synchronized = call_black_white & (~vsync);
        call_edge_detection_synchronized = call_edge_detection & (~vsync);
    end

    // BW entity: black_white (actually grey) filter; reads from buf1 and writes into buf1
    do_black_white do_black_white_inst(
        .rst_i(reset_BW_entity),
        .clk_i(clk_25_vga),
        .enable_filter(call_black_white_synchronized),
        .led_done(done_BW_from_module),
        .rdaddr_buf1(rdaddress_buf1_from_do_BW), // goes to mux of rdaddress_buf_1
        .din_buf1(rddata_buf_1), // comes from out of buf1
        .wraddr_buf1(wraddress_buf1_from_do_BW), // goes to mux of wraddress_buf_2
        .dout_buf1(wrdata_buf1_from_do_BW), // goes to mux of wrdata_buf_2
        .we_buf1(wren_buf1_from_do_BW) // goes to mux of wren_buf_2
    );

    // ED entity: Sobel edge detection; reads from buf2 and writes into buf2
    do_edge_detection do_edge_detection_inst(
        .rst_i(reset_ED_entity),
        .clk_i(clk_25_vga),
        .enable_sobel_filter(call_edge_detection_synchronized),
        .led_sobel_done(done_ED_from_module),
        .rdaddr_buf1(rdaddress_buf1_from_do_ED), // goes to mux of rdaddress_buf_1
        .din_buf1(rddata_buf_1), // comes from out of buf1
        .wraddr_buf2(wraddress_buf2_from_do_ED), // goes to mux of wraddress_buf_2
        .dout_buf2(wrdata_buf2_from_do_ED), // goes to mux of wrdata_buf_2
        .we_buf2(wren_buf2_from_do_ED) // goes to mux of wren_buf_2
    );

endmodule
